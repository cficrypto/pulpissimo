// BACCTODO verify that this does not interfere with parameters
`ifndef CFI_INSTR_WIDTH_DEF
`define CFI_INSTR_WIDTH_DEF 40
`endif